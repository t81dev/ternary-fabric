/*
 * Vector Engine: TFM-Compliant Parallel Ternary Processor
 * Tiles 'N' Ternary Processing Elements (TPEs) for SIMD operations.
 * Implements Logical Mapping: Offset = (depth * LANES) + lane_id
 */
module vector_engine #(
    parameter LANES = 16,           // Configurable SIMD width
    parameter ACCUM_WIDTH = 32      // Binary precision per lane
)(
    input  wire                     clk,
    input  wire                     reset,
    
    // Control Interface
    input  wire                     enable,
    input  wire [2:0]               op_mode,      // Command: 01=Dot, etc.
    
    // Data Interface (Unpacked from PT-5 by upstream Bus Controller)
    input  wire [(LANES*2)-1:0]     bus_weights,  // 2-bits per lane
    input  wire [(LANES*2)-1:0]     bus_inputs,   // 2-bits per lane
    
    // Output: Parallel Accumulator State
    output wire [(LANES*ACCUM_WIDTH)-1:0] vector_out
);

    genvar i;
    generate
        for (i = 0; i < LANES; i = i + 1) begin : gen_lanes
            // Instantiate the TPE for each lane
            ternary_lane_alu lane_inst (
                .clk(clk),
                .reset(reset),
                .enable(enable),
                .op_mode(op_mode),        // <--- FIXED: Passing the command down
                .weight(bus_weights[i*2 +: 2]),
                .trit_in(bus_inputs[i*2 +: 2]),
                .accumulator(vector_out[i*ACCUM_WIDTH +: ACCUM_WIDTH])
            );
        end
    endgenerate

endmodule